// soc_system.v

// Generated using ACDS version 13.1 162 at 2019.01.02.20:41:33

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        reset_reset_n,                           //                       reset.reset_n
		output wire [14:0] memory_mem_a,                            //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                           //                            .mem_ba
		output wire        memory_mem_ck,                           //                            .mem_ck
		output wire        memory_mem_ck_n,                         //                            .mem_ck_n
		output wire        memory_mem_cke,                          //                            .mem_cke
		output wire        memory_mem_cs_n,                         //                            .mem_cs_n
		output wire        memory_mem_ras_n,                        //                            .mem_ras_n
		output wire        memory_mem_cas_n,                        //                            .mem_cas_n
		output wire        memory_mem_we_n,                         //                            .mem_we_n
		output wire        memory_mem_reset_n,                      //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                           //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                          //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                        //                            .mem_dqs_n
		output wire        memory_mem_odt,                          //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                           //                            .mem_dm
		input  wire        memory_oct_rzqin,                        //                            .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,         //                      hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,           //                            .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,           //                            .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,           //                            .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,           //                            .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,           //                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,           //                            .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,            //                            .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,         //                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,         //                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,         //                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,           //                            .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,           //                            .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,           //                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,             //                            .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,             //                            .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,             //                            .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,             //                            .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,             //                            .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,             //                            .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,             //                            .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,              //                            .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,              //                            .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,             //                            .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,              //                            .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,              //                            .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,              //                            .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,              //                            .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,              //                            .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,              //                            .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,              //                            .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,              //                            .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,              //                            .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,              //                            .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,             //                            .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,             //                            .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,             //                            .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,             //                            .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,            //                            .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,           //                            .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,           //                            .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,            //                            .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,             //                            .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,             //                            .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,             //                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,             //                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,             //                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,             //                            .hps_io_i2c1_inst_SCL
		output wire        hps_h2f_reset_reset_n,                   //               hps_h2f_reset.reset_n
		input  wire        clk_clk,                                 //                         clk.clk
		output wire        hps_terminal_conduit_end_main_reset_n,   //    hps_terminal_conduit_end.main_reset_n
		output wire        hps_terminal_conduit_end_rd,             //                            .rd
		input  wire        hps_terminal_conduit_end_rd_valid,       //                            .rd_valid
		input  wire [63:0] hps_terminal_conduit_end_rd_instruction, //                            .rd_instruction
		output wire        hps_terminal_conduit_end_wr,             //                            .wr
		input  wire        hps_terminal_conduit_end_wr_busy,        //                            .wr_busy
		output wire [63:0] hps_terminal_conduit_end_wr_instruction, //                            .wr_instruction
		output wire [31:0] pio_led_external_connection_export       // pio_led_external_connection.export
	);

	wire  [31:0] mm_interconnect_0_hps_terminal_avalon_slave_writedata; // mm_interconnect_0:HPS_Terminal_avalon_slave_writedata -> HPS_Terminal:s_writedata
	wire   [9:0] mm_interconnect_0_hps_terminal_avalon_slave_address;   // mm_interconnect_0:HPS_Terminal_avalon_slave_address -> HPS_Terminal:s_address
	wire         mm_interconnect_0_hps_terminal_avalon_slave_write;     // mm_interconnect_0:HPS_Terminal_avalon_slave_write -> HPS_Terminal:s_write
	wire         mm_interconnect_0_hps_terminal_avalon_slave_read;      // mm_interconnect_0:HPS_Terminal_avalon_slave_read -> HPS_Terminal:s_read
	wire  [31:0] mm_interconnect_0_hps_terminal_avalon_slave_readdata;  // HPS_Terminal:s_readdata -> mm_interconnect_0:HPS_Terminal_avalon_slave_readdata
	wire         hps_h2f_axi_master_awvalid;                            // hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	wire   [2:0] hps_h2f_axi_master_arsize;                             // hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	wire   [1:0] hps_h2f_axi_master_arlock;                             // hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	wire   [3:0] hps_h2f_axi_master_awcache;                            // hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	wire         hps_h2f_axi_master_arready;                            // mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	wire  [11:0] hps_h2f_axi_master_arid;                               // hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	wire         hps_h2f_axi_master_rready;                             // hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	wire         hps_h2f_axi_master_bready;                             // hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	wire   [2:0] hps_h2f_axi_master_awsize;                             // hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	wire   [2:0] hps_h2f_axi_master_awprot;                             // hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	wire         hps_h2f_axi_master_arvalid;                            // hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	wire   [2:0] hps_h2f_axi_master_arprot;                             // hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	wire  [11:0] hps_h2f_axi_master_bid;                                // mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	wire   [3:0] hps_h2f_axi_master_arlen;                              // hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	wire         hps_h2f_axi_master_awready;                            // mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	wire  [11:0] hps_h2f_axi_master_awid;                               // hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	wire         hps_h2f_axi_master_bvalid;                             // mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	wire  [11:0] hps_h2f_axi_master_wid;                                // hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	wire   [1:0] hps_h2f_axi_master_awlock;                             // hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	wire   [1:0] hps_h2f_axi_master_awburst;                            // hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	wire   [1:0] hps_h2f_axi_master_bresp;                              // mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	wire   [3:0] hps_h2f_axi_master_wstrb;                              // hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	wire         hps_h2f_axi_master_rvalid;                             // mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	wire  [31:0] hps_h2f_axi_master_wdata;                              // hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	wire         hps_h2f_axi_master_wready;                             // mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	wire   [1:0] hps_h2f_axi_master_arburst;                            // hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	wire  [31:0] hps_h2f_axi_master_rdata;                              // mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	wire  [29:0] hps_h2f_axi_master_araddr;                             // hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	wire   [3:0] hps_h2f_axi_master_arcache;                            // hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	wire   [3:0] hps_h2f_axi_master_awlen;                              // hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	wire  [29:0] hps_h2f_axi_master_awaddr;                             // hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	wire  [11:0] hps_h2f_axi_master_rid;                                // mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	wire         hps_h2f_axi_master_wvalid;                             // hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	wire   [1:0] hps_h2f_axi_master_rresp;                              // mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	wire         hps_h2f_axi_master_wlast;                              // hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	wire         hps_h2f_axi_master_rlast;                              // mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                  // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;               // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire         mm_interconnect_0_pio_led_s1_write;                    // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                 // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;         // mm_interconnect_0:sysID_control_slave_address -> sysID:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;        // sysID:readdata -> mm_interconnect_0:sysID_control_slave_readdata
	wire  [31:0] hps_f2h_irq0_irq;                                      // irq_mapper:sender_irq -> hps:f2h_irq_p0
	wire  [31:0] hps_f2h_irq1_irq;                                      // irq_mapper_001:sender_irq -> hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [HPS_Terminal:s_reset, mm_interconnect_0:sysID_reset_reset_bridge_in_reset_reset, pio_led:reset_n, sysID:reset_n]
	wire         rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	soc_system_hps #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.h2f_rst_n                (hps_h2f_reset_reset_n),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_h2f_axi_master_awid),         //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_h2f_axi_master_awaddr),       //                  .awaddr
		.h2f_AWLEN                (hps_h2f_axi_master_awlen),        //                  .awlen
		.h2f_AWSIZE               (hps_h2f_axi_master_awsize),       //                  .awsize
		.h2f_AWBURST              (hps_h2f_axi_master_awburst),      //                  .awburst
		.h2f_AWLOCK               (hps_h2f_axi_master_awlock),       //                  .awlock
		.h2f_AWCACHE              (hps_h2f_axi_master_awcache),      //                  .awcache
		.h2f_AWPROT               (hps_h2f_axi_master_awprot),       //                  .awprot
		.h2f_AWVALID              (hps_h2f_axi_master_awvalid),      //                  .awvalid
		.h2f_AWREADY              (hps_h2f_axi_master_awready),      //                  .awready
		.h2f_WID                  (hps_h2f_axi_master_wid),          //                  .wid
		.h2f_WDATA                (hps_h2f_axi_master_wdata),        //                  .wdata
		.h2f_WSTRB                (hps_h2f_axi_master_wstrb),        //                  .wstrb
		.h2f_WLAST                (hps_h2f_axi_master_wlast),        //                  .wlast
		.h2f_WVALID               (hps_h2f_axi_master_wvalid),       //                  .wvalid
		.h2f_WREADY               (hps_h2f_axi_master_wready),       //                  .wready
		.h2f_BID                  (hps_h2f_axi_master_bid),          //                  .bid
		.h2f_BRESP                (hps_h2f_axi_master_bresp),        //                  .bresp
		.h2f_BVALID               (hps_h2f_axi_master_bvalid),       //                  .bvalid
		.h2f_BREADY               (hps_h2f_axi_master_bready),       //                  .bready
		.h2f_ARID                 (hps_h2f_axi_master_arid),         //                  .arid
		.h2f_ARADDR               (hps_h2f_axi_master_araddr),       //                  .araddr
		.h2f_ARLEN                (hps_h2f_axi_master_arlen),        //                  .arlen
		.h2f_ARSIZE               (hps_h2f_axi_master_arsize),       //                  .arsize
		.h2f_ARBURST              (hps_h2f_axi_master_arburst),      //                  .arburst
		.h2f_ARLOCK               (hps_h2f_axi_master_arlock),       //                  .arlock
		.h2f_ARCACHE              (hps_h2f_axi_master_arcache),      //                  .arcache
		.h2f_ARPROT               (hps_h2f_axi_master_arprot),       //                  .arprot
		.h2f_ARVALID              (hps_h2f_axi_master_arvalid),      //                  .arvalid
		.h2f_ARREADY              (hps_h2f_axi_master_arready),      //                  .arready
		.h2f_RID                  (hps_h2f_axi_master_rid),          //                  .rid
		.h2f_RDATA                (hps_h2f_axi_master_rdata),        //                  .rdata
		.h2f_RRESP                (hps_h2f_axi_master_rresp),        //                  .rresp
		.h2f_RLAST                (hps_h2f_axi_master_rlast),        //                  .rlast
		.h2f_RVALID               (hps_h2f_axi_master_rvalid),       //                  .rvalid
		.h2f_RREADY               (hps_h2f_axi_master_rready),       //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (),                                // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (),                                //                  .awaddr
		.h2f_lw_AWLEN             (),                                //                  .awlen
		.h2f_lw_AWSIZE            (),                                //                  .awsize
		.h2f_lw_AWBURST           (),                                //                  .awburst
		.h2f_lw_AWLOCK            (),                                //                  .awlock
		.h2f_lw_AWCACHE           (),                                //                  .awcache
		.h2f_lw_AWPROT            (),                                //                  .awprot
		.h2f_lw_AWVALID           (),                                //                  .awvalid
		.h2f_lw_AWREADY           (),                                //                  .awready
		.h2f_lw_WID               (),                                //                  .wid
		.h2f_lw_WDATA             (),                                //                  .wdata
		.h2f_lw_WSTRB             (),                                //                  .wstrb
		.h2f_lw_WLAST             (),                                //                  .wlast
		.h2f_lw_WVALID            (),                                //                  .wvalid
		.h2f_lw_WREADY            (),                                //                  .wready
		.h2f_lw_BID               (),                                //                  .bid
		.h2f_lw_BRESP             (),                                //                  .bresp
		.h2f_lw_BVALID            (),                                //                  .bvalid
		.h2f_lw_BREADY            (),                                //                  .bready
		.h2f_lw_ARID              (),                                //                  .arid
		.h2f_lw_ARADDR            (),                                //                  .araddr
		.h2f_lw_ARLEN             (),                                //                  .arlen
		.h2f_lw_ARSIZE            (),                                //                  .arsize
		.h2f_lw_ARBURST           (),                                //                  .arburst
		.h2f_lw_ARLOCK            (),                                //                  .arlock
		.h2f_lw_ARCACHE           (),                                //                  .arcache
		.h2f_lw_ARPROT            (),                                //                  .arprot
		.h2f_lw_ARVALID           (),                                //                  .arvalid
		.h2f_lw_ARREADY           (),                                //                  .arready
		.h2f_lw_RID               (),                                //                  .rid
		.h2f_lw_RDATA             (),                                //                  .rdata
		.h2f_lw_RRESP             (),                                //                  .rresp
		.h2f_lw_RLAST             (),                                //                  .rlast
		.h2f_lw_RVALID            (),                                //                  .rvalid
		.h2f_lw_RREADY            (),                                //                  .rready
		.f2h_irq_p0               (hps_f2h_irq0_irq),                //          f2h_irq0.irq
		.f2h_irq_p1               (hps_f2h_irq1_irq)                 //          f2h_irq1.irq
	);

	soc_system_sysID sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	HPS_Terminal hps_terminal (
		.s_clk          (clk_clk),                                               //   clock_sink.clk
		.s_reset        (rst_controller_reset_out_reset),                        //   reset_sink.reset
		.s_write        (mm_interconnect_0_hps_terminal_avalon_slave_write),     // avalon_slave.write
		.s_read         (mm_interconnect_0_hps_terminal_avalon_slave_read),      //             .read
		.s_address      (mm_interconnect_0_hps_terminal_avalon_slave_address),   //             .address
		.s_writedata    (mm_interconnect_0_hps_terminal_avalon_slave_writedata), //             .writedata
		.s_readdata     (mm_interconnect_0_hps_terminal_avalon_slave_readdata),  //             .readdata
		.main_reset_n   (hps_terminal_conduit_end_main_reset_n),                 //  conduit_end.export
		.rd             (hps_terminal_conduit_end_rd),                           //             .export
		.rd_valid       (hps_terminal_conduit_end_rd_valid),                     //             .export
		.rd_instruction (hps_terminal_conduit_end_rd_instruction),               //             .export
		.wr             (hps_terminal_conduit_end_wr),                           //             .export
		.wr_busy        (hps_terminal_conduit_end_wr_busy),                      //             .export
		.wr_instruction (hps_terminal_conduit_end_wr_instruction)                //             .export
	);

	soc_system_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_h2f_axi_master_awid                                        (hps_h2f_axi_master_awid),                               //                                       hps_h2f_axi_master.awid
		.hps_h2f_axi_master_awaddr                                      (hps_h2f_axi_master_awaddr),                             //                                                         .awaddr
		.hps_h2f_axi_master_awlen                                       (hps_h2f_axi_master_awlen),                              //                                                         .awlen
		.hps_h2f_axi_master_awsize                                      (hps_h2f_axi_master_awsize),                             //                                                         .awsize
		.hps_h2f_axi_master_awburst                                     (hps_h2f_axi_master_awburst),                            //                                                         .awburst
		.hps_h2f_axi_master_awlock                                      (hps_h2f_axi_master_awlock),                             //                                                         .awlock
		.hps_h2f_axi_master_awcache                                     (hps_h2f_axi_master_awcache),                            //                                                         .awcache
		.hps_h2f_axi_master_awprot                                      (hps_h2f_axi_master_awprot),                             //                                                         .awprot
		.hps_h2f_axi_master_awvalid                                     (hps_h2f_axi_master_awvalid),                            //                                                         .awvalid
		.hps_h2f_axi_master_awready                                     (hps_h2f_axi_master_awready),                            //                                                         .awready
		.hps_h2f_axi_master_wid                                         (hps_h2f_axi_master_wid),                                //                                                         .wid
		.hps_h2f_axi_master_wdata                                       (hps_h2f_axi_master_wdata),                              //                                                         .wdata
		.hps_h2f_axi_master_wstrb                                       (hps_h2f_axi_master_wstrb),                              //                                                         .wstrb
		.hps_h2f_axi_master_wlast                                       (hps_h2f_axi_master_wlast),                              //                                                         .wlast
		.hps_h2f_axi_master_wvalid                                      (hps_h2f_axi_master_wvalid),                             //                                                         .wvalid
		.hps_h2f_axi_master_wready                                      (hps_h2f_axi_master_wready),                             //                                                         .wready
		.hps_h2f_axi_master_bid                                         (hps_h2f_axi_master_bid),                                //                                                         .bid
		.hps_h2f_axi_master_bresp                                       (hps_h2f_axi_master_bresp),                              //                                                         .bresp
		.hps_h2f_axi_master_bvalid                                      (hps_h2f_axi_master_bvalid),                             //                                                         .bvalid
		.hps_h2f_axi_master_bready                                      (hps_h2f_axi_master_bready),                             //                                                         .bready
		.hps_h2f_axi_master_arid                                        (hps_h2f_axi_master_arid),                               //                                                         .arid
		.hps_h2f_axi_master_araddr                                      (hps_h2f_axi_master_araddr),                             //                                                         .araddr
		.hps_h2f_axi_master_arlen                                       (hps_h2f_axi_master_arlen),                              //                                                         .arlen
		.hps_h2f_axi_master_arsize                                      (hps_h2f_axi_master_arsize),                             //                                                         .arsize
		.hps_h2f_axi_master_arburst                                     (hps_h2f_axi_master_arburst),                            //                                                         .arburst
		.hps_h2f_axi_master_arlock                                      (hps_h2f_axi_master_arlock),                             //                                                         .arlock
		.hps_h2f_axi_master_arcache                                     (hps_h2f_axi_master_arcache),                            //                                                         .arcache
		.hps_h2f_axi_master_arprot                                      (hps_h2f_axi_master_arprot),                             //                                                         .arprot
		.hps_h2f_axi_master_arvalid                                     (hps_h2f_axi_master_arvalid),                            //                                                         .arvalid
		.hps_h2f_axi_master_arready                                     (hps_h2f_axi_master_arready),                            //                                                         .arready
		.hps_h2f_axi_master_rid                                         (hps_h2f_axi_master_rid),                                //                                                         .rid
		.hps_h2f_axi_master_rdata                                       (hps_h2f_axi_master_rdata),                              //                                                         .rdata
		.hps_h2f_axi_master_rresp                                       (hps_h2f_axi_master_rresp),                              //                                                         .rresp
		.hps_h2f_axi_master_rlast                                       (hps_h2f_axi_master_rlast),                              //                                                         .rlast
		.hps_h2f_axi_master_rvalid                                      (hps_h2f_axi_master_rvalid),                             //                                                         .rvalid
		.hps_h2f_axi_master_rready                                      (hps_h2f_axi_master_rready),                             //                                                         .rready
		.clk_clk_clk                                                    (clk_clk),                                               //                                                  clk_clk.clk
		.hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysID_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                        //                        sysID_reset_reset_bridge_in_reset.reset
		.HPS_Terminal_avalon_slave_address                              (mm_interconnect_0_hps_terminal_avalon_slave_address),   //                                HPS_Terminal_avalon_slave.address
		.HPS_Terminal_avalon_slave_write                                (mm_interconnect_0_hps_terminal_avalon_slave_write),     //                                                         .write
		.HPS_Terminal_avalon_slave_read                                 (mm_interconnect_0_hps_terminal_avalon_slave_read),      //                                                         .read
		.HPS_Terminal_avalon_slave_readdata                             (mm_interconnect_0_hps_terminal_avalon_slave_readdata),  //                                                         .readdata
		.HPS_Terminal_avalon_slave_writedata                            (mm_interconnect_0_hps_terminal_avalon_slave_writedata), //                                                         .writedata
		.pio_led_s1_address                                             (mm_interconnect_0_pio_led_s1_address),                  //                                               pio_led_s1.address
		.pio_led_s1_write                                               (mm_interconnect_0_pio_led_s1_write),                    //                                                         .write
		.pio_led_s1_readdata                                            (mm_interconnect_0_pio_led_s1_readdata),                 //                                                         .readdata
		.pio_led_s1_writedata                                           (mm_interconnect_0_pio_led_s1_writedata),                //                                                         .writedata
		.pio_led_s1_chipselect                                          (mm_interconnect_0_pio_led_s1_chipselect),               //                                                         .chipselect
		.sysID_control_slave_address                                    (mm_interconnect_0_sysid_control_slave_address),         //                                      sysID_control_slave.address
		.sysID_control_slave_readdata                                   (mm_interconnect_0_sysid_control_slave_readdata)         //                                                         .readdata
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                 //       clk.clk
		.reset      (),                 // clk_reset.reset
		.sender_irq (hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset_n),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
