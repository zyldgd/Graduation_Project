��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e��T`U���kO_:��(R��]͋�}�X`ׂ��O��Х)\������}r�����x T�Q.��ב{�@g��^�Q�S��t�Ds� z{3aT�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���	e��"a5���f���wR����.F�o!��5���?��Ԣ*5lkc�Bڝ������t�}�8���Ok�>�ځJ"�ꄢݬ�"4'4����^�0L����܃��x ~b��4�b��@��E"�Fu��(���f������~X�2S!���r�E/�=�A��G'ş��6�J�Y��,�bd�C�S��ٌ0�{Jؖ����E���͚�<۳�7�;�@k�ރ͍�B~R���,��^u��\@������DWa�!�Tָ�L���%��V�9���*�e���c� ґ1��rLmo�B�jV��F�7Rݖ�����}���݌DkJGh����!��|,��*zjf�p�Q�DǕ�Q�C�#�{=F�9������E��R@k���>v�����"�S��"��[`v��U�7�� J��O�nC�$d�D�a|o�P���e�=?�D�Q�	���D���<x��dڴtRy��bO�I�� @�a�����a�Wy��'�_�����Y�7�ߦ��f0�}Q���'
���X�[l��hm��UA�x���ك甒t�G�G���i|Y�ot��\��5��8�������SLm��.�pJf��:5F0zOw�����bD.�0�N7ɘ/�K5���s�ߛ&���ǡ	��P ��s����/���|+gj��/�&�Edi(K$>6v��w�co@ҍki�X?����	E��*�)���ʴ�SѱZ�-�7+��so�k���=��|�M.�2�m�2��[^�[p�>s�l���-����)b}jD��ܗ�'h�����+-�HH&�jH`��x�U3Ԍ�R�`�$��)����#n��	��_�\!��k]�'V�r�p�p��91���	��w3?i�)D6/!&V�1�v�B�Q�G-���_H�$�3sT2K�jC�\�˦�6`��󁷴�P�ј���E :�7,�dmY��ދ�g.��p�R�޹q�6��>�U�����x�0��z�l�h|���3�=��\q�x�u!�X�V��)�	��g0����[{+��#ԟg�g�?'Y"=�{dg��<��q�հ���y���v$3�Y�nO�1E��ra�@����<ZhU��İ[�ms��_7E�!c7J�E����џ�^�̍|���$t�ZM�������(%	���(Ib4F���G�ߒ�I%�����$���X����ҺS��)6C����WDs6,�>��ʽ�c���'��T�QJ0ة�`����-�R �yr|b9���	T׀�xΜ��A���cto�}��t�a��kq3�(_�ȼN�A�5O�.�_���!��,���B�@��;H0
�;��2�]Y�6�Ԃ�ih�Xe��u�<���$�P��jl�ם�[���z%4�'���0�
�[�v�Ĕ��(m[z�S"���^�ϹI�B�J��'�x.=�ei�,V��m��W��b>�(�_+ʧ�"]>����ޖ<]�1�ز��[��K�����P���*�|��;��j������B�l����mX�0��{������cW�[�R��}���Z��xwnm�t���d�Z �f-�~������>���R�!^�;��qq飘��\�
���}&��������+�.�A�1�M��w*���72H�A��1xxw��%�V���S5���z�J��Wզ���ʨ5���;Xh�>�a�h~����	Y�3����#t8�G�������*wcU���w��W�;'����&�0�"���.�_���u��,��%�� ���p��Z�q�~Y��	��T�(p2���6o��̊�G!K���1���)dX��0(���B���@�}�Cl�}��� ���߭R�Ր�biI���?}���#��XN�qS>�H�`L��˞6$ ���<O�L]�0�/�83q� \�q�+��K渄˯����0(�n�ŷ����CO(�^�1pgM"����p���r��6�~{^�Ep]��4��c0��<��4�#�o��%�b�^Q��8�F��{�>��U[1_�2��*8O�.��hg���@�Q![b�E|꣥���_��a��tM��g���� ��l� q���\�!X�p��S; �����#�5^���č���I�GaBAU8���d�S#�&�E�m�7�(�vN��
4�v�|��S�nK��P�Z72;�N?�V�O�����d�M%��]@F�E�\f$�t�ĵ����aw�_��6IlZx
��JP�eje$��?|��ﱣ&�]:��}F���=�e���$��fR�U��.ޫ`���Oa��>p�����9�}�Z� v���0��$("�q����V��k��k��ě��6��	�_��O����ƙ����wo�����L�oE�9����~i}��S�B)X F�v��˜��m�� U� �ʱ��p����
���#/�5ADj�D5����l�����\)�ZI�8E��g�ᴚG;Z����.��H肯�-7�����X�b��.� ���MC�1�9όYE��	A�����Z�U�t0�N^lF�!�<W�ʻ+!�����50�\�K�j��5�%�)��Z�77���z���2������߆s��L1��0H�1ɺ)��O{<����� /9̲Z��[���S�2�T؎����/�E@���N9-�u%�MȤ�"��
��(I�25j�ڔ(o��Fz�7��,�2Їzq��_�F�� �O��V{��r��t��1���d����(Qk�[��Ю��N��$)�s�ѷ$!�p�8�gg���w��u����k�(�:v����'N	�&�?'oXX*�n(o��&JR[�KA�ۮ3��8�!��{��f�\� �M�>΁~�Ч�{1m�d�7֔�1�����^3?��vv�!ؕ��#�`�M�,�
Q4��d�vY �c��M�y�J�n���GC�p��#y��fF��6�-�S��+��YpV�JY7K�)٧�͗MG��%�怖'�e�B�2`w9:�P�BbQ�����1��Y�^�� e�a�N�J� �Y���o�Ơ��G|m������o��/�l ��c���Lr�:���7J3�$D_4�Y�#����[��]h�W~]6��@L����x�m|$P�.I!Y7�L���F�b�5HV����n��|c�U_�$<��J�!m|�����m���1�_Z��`u�d驗�A��Vxh=DZ��q_�NH�%�Ij�-m��(yQ�ޟ?�r���6��`�"�_�Z}r�0*_� $g��>]G�??�)���(f@jlZ�E�19�j݅�@������\3�T�8SJ�#Q9�l 67~�)�:����&"Ǡ����� �BG����\Hڪ&.�ˡ� ]Ie�aL�.zZ�^#م��υ:�D�v��Y��nOS�}�R�cǐ4=��^r��&{�ܻ�5�����.ۼ%Sw���(i�B>U�CU�O��ߔ���k��xk��9�ܢr�+���G�^U
��A�� η�H��z��/�7�*a|�0P�/o�E��I�ߎ9�$7�:y,
���-!i���p���%DՋ"*�f�8�Y�>
ῐ�Ѵ��+��6�ͭ��D2:{\,0=+�T��i^YD���=Ӳ�F�O:e�a��h#�w�(���Gܼ�Xkc�8,_J�������0� 4H�<���#�)���Ϝ��?I	��>Ԇg-s��0:��VYh�
�Y�qք�ur����Eh
Q�A�����ć,���d�i��ǏM����!���>�E��}�#�sѐ�s� ;��V ��t{��28�ڈ�m�,>�rwW�C�e�Vaξ�����S�2� r��c���m�,�ʿ�GU5��x{t�=��uG�p���E�ы@��p�
f���gqep���<�
�#���oҶ�	�H�2�P�+�:���d 1��h��� ��@k"Ş�S�,��q�c�IX�\AF]�}��d�3՘�Ӳ�wdn�Y?5%n�Z�Y�}y��Gm�Ld����F�\mQ5;�� ��S��Xt��v��F�V�Jn��'V.$Yل�`*���N�w�ht��:8�Ҳ2{e��]��Yv˵���k��$�Z ,-�xiG��}2�6K|h�5w#>PK���e'�D"[w�
{�5��벦���MF�:�K�3W�>Z�B��������P�Vpv��q	C������ӯ*�D���qy��H(�R\��U�����V"����rԓ�V�ֆ��vn@�A�A��u�- �R���l0�����z�5����ɯd�R[&u���b�]�K�k%�De���A!Bl�+�����w0����� �Av׃�g���$X��dyf�w~����5���ꥢ�~H��a�ۘ�5�	���%�#M)[����#�C�a�,<��%��<_0�jG�;qے���3��ù;��G2�R��^�=b�iR;c�-ÑOq
Z��������1������ş�����XH<�����o�P�E%��sms���u��j,
%-�m�xǯ�f�UI��\.I ��,��n�%�7�-
��R��X�ƨ����J�q!���ﾻzKf/��Ѷ���Cp^��^U{焸F�z]Ao����Z����8��#v��R�T5�#α��_�����T�~!�  8��
̿��-[M���8l�����n��@�7�T U�x3������ؑo���f�7��W#�����pA:��R<�@��� z��U�I�FM�� (�'��ǯ�I�P%3)@�i�!�g���La$)�N��"��}n�tCP�5�]^a�Y��{V���O0B�_`�C_){O��o�������~I���ݼRۈ�x�ڵ���o�Uv��5��ȯ�����Dٜ%Z絋�ԁL����v����|����1�� e�|�)���|{�W�k�z��¼''����p�-}��
���I�o(�uK1���3:6�JtCjBr�D����Z��b	�
�S�T��vG��ݷu�jAm��!m�i��@+�M�)��y��/o`(uqV���R�%͞���(TJ�D��sr����\����C�*���&�A54[���͜6v:Jj�U��/Ԗ�Y[$�;nwk��nM>�n+�¼z�㘪�أҗ!�m�0ٯ�� ��:���M9Zͳkru4}P>0�	�6�)c����gc�>e�v�Y42%P���"w�E�*ڒ6a�G�hz*�qɜ���>�>��:� �
HS�-���a�
ge�C���=�$�q�`ߘ�q��K0,)r�4�G�G}g�N����֎=����e�?����굒"Ɂ)�1�z�)mG�Ew{^��,:��6��vu�����3���S�v���&\vwu
+�*�6G��g#�e���	wf�o%Ϡ�^��u;��w����jj��]��A����J�(�L���,&Lm����qs��m����0~a�`���*Y����"��M������M�+N�Y�u���Ē%�f��6>�=��s��AAu�H%%�> �Th,@���tQL�@�'�.�������F|*�0ħ��|��lF�ti˩V ��P�y����ť
r��fp���V�v�����7e����2`?�ӎ?��ir�f��fh94�	7�N� ��5����X�q�Mr:�/���b�\r	t��.�� �8��s�o�~W�r"���P^�ݤ�w��Hl�,����*
x�i�����(H� �}�';��FL)Ͼ��'��i�4+��3
�Ʋv�'d]��]��ca^vR9�<o�YW��OAo�b�&�7�]y<���I��ʮt:�rEE���]�BDm~s�{�d,��v�ٷjQ�G�Ĺ��D�b�LR�ջ1C�B� )�s0��
.:=����k���sb�l��H��ֲ��=�V>{���?	\��v�7;����n��.��ԔZ������F ��y��5�G���n�Ӻ���7��p�Z��>���?����R���S�S12��}���|�xI��~��1�&@c[���3�t���߀�q�A�@4�!0�'��k�����4���dr�r$�J�&������A9pu�_�X��#��.�)���h0����Ћ����,��b�;�ԇ<^&�e9��u,X�U�I/�hV ��NU�3��nr*��n>}��{.�e�Tg�<%95kL�����ki�_ug�K�1�3A2.ȴ����|�N��Ʒ�V1�����9=<�0Wiသ�S�"$�ŎD��T�_6��H�� F6�b=�VD]}�X|��kad��8n��ª�T��=�0���1���s}����R�N/���?���[A���s�vP���QP�S�X����d��;S��Y�C������!öv�� X	wY�D�of�YN��I��K�&y��{)�;]�Ʒ��ESY��_}�=p�3LwUi��;�	��y���7�ԙ�����7�Ц�`�b���Οy]�x�ؙ�&d��$#i�����?�x ��(rD�8Uw�_��U�%m�iezx�dl(ò�gM�w�E���%�,vگ�l���r�b�����U��K�����&RZe5H?=G���j9��� ˋ��U��r5*.��h��H��+��W��nZ~ᢵ�&�o�vSw��#v�ǭH&b�c����Um���=X>��mh�-�vl�������f��~�y5F��N�{����gy��	��st�I�Xl�ei�n�TC�� }��jZTu���Ϥ�N�2�v���gՅj�?��[p�ܐ����O@��@J����D�:@�禍W&\ :!��I<�U����K�_�S��
ѩ�>��_�@X?;_
�g�k[l����5��\�͑l�Ԭ�#ऒ�7�usG��hB	{�}�>'1e�I���_��|��_9.��!��?��S�����Y�;�8�H��5�=wT��;����m}4g�I{rz|q���t'D��}�������>ic���btnm!�"E�G8%�޴�y~�>	�[ދ��h���D&KK	�o�`I	��%��Ũ�v�j@(%�G�W�z:{��x�f&p_Mw����p»mKGr`��b�I�Ʃs^}�gJ1޷��6$�_K.X�*�[-c�f;�p�[���-�	���ά[/���6)ğI�͢\��.��z�&dD� �kNg���h��Դu�	�&�!�o:��\SىL�'�️�_挣�֕���]����8�:$g�;����65�n�xڐC�0�4
�*����˱L��9�'��,��25�4�o�V��A6	}�k�	VƆѓ��N��!A�)�'; N�#6�����{~P]'l
K�XU(k?(�ʰ�8K{o�|@��ˆ
l_Y�.	h��m XF眖DJ�f�J&�6{�J��'Ep"�$����<A7���jH�\	 �gx�pp9����ln��Z#m{�v>�BE�l�"�ݮ�{�|+��
B"៑N�r>�/B��Xj��I�7�sDR#��L���K���n�!P���4f2c#�9�F��z�gl�;�Ix��RCK���;p�uz��D�r��_�G�j�
w8��dAv��·��R+Y2$����!���"�T��"�����J�8�C0��R-�Xj�_9E/q��!�(2��by�rn�#��/�ɍ�}�X��&e5���p���^*�0�]�/�(d}��N�5uA���بy*����7qJ���?�/�AMO�Y��W�EH�M��bB��i��}H:�L����T���>���L}����3�0��E;��'�ҕ�2�*T9
~��Wg9vL���cS���D?��������0l���0$y�G��N���JvOg�a� TŌ��^ PO|t�v��g�Qv�t��k%�%M�s���ڏ^@��A�x��D"�����^:�w��p�E_� �ͱ���HӽmK2%]�۬84�Uw�D����z��H&D6��w!����W���X�n���[Fa�M&�n�+����Q�gk���$�Ï�=+ː�S tM�wE<�lF⻩���b�7��H�D�r�68��T���v�݌���CbK:s����w߼1#32<�'�Ѥ�[�c���y��v���(o��kS�i�S�ioϠ����j5�ʗڇ�K.����<�k�q?)3P����[�1��1~y��j���3Ԣ���ܙ�
�8��j{�X�j@�^�%�aM��Fev�i��$]�^r�,��>�ePG,B��\�P��gk�L��"��R�A�f�)�����P��Vi�k���,r,��>s���4�Ł�L�R ��i�A��10ܥ���&1����XA��|����1�n�y�)�!��B>2`�C�ċ��'�L��s�p3��N[8����?�,���,��Mu {�R��B���?v��دx���X Z=t?���[{g�[8�V��&I�l!��~��F��\�Q �� Sg��@@�4�F�!)��a�U4r��ڴ.�n�g5��mY���^�{�6F��B��޾����c���XW+u���Ɩ�gK�����ǀ�f�(�:4F+� h7Vy�S]lni�k���ug�}�+##���(B�I�-[�4S΋A?��ژg�X��%�2C>�f�UN�~�5�lOm��<]�dl8#�j��gg�-�ѣ/�?V�&lx��AXPQ��Y�P*����IvxhJޜ9���vz`��ˮ���ш7ɍ��e��Dk��K�@$cUfI�\�C������{�C�����k��p�y�
�HnL�7�,S�]�[I�ѣ��-N,b[��Y�C^��|�g� ��@Y���R�j�,������<���W�!�����
�\N��a^�3��-5�>���-.%�՚T��ʃ��[r�8Z��G����R�h1
u�����>�'-9uB�Aq�����e٤��[XC��]M^� �/�O>!�X��)M��oĘ���G������äm̮?o�5Z���ͦp���.M̰8 ol�8"9���(�}��H���*���G�����c�v:���%�^w���$�u�ق�s�mnL�Z�� �@�ڏ��'D�(z�8@���S�L@1]g�����dqLj$�(���ڱ�3��΂'����hin�8�r�Ȱ�N }Na&=N3��`6;B��	�����P	�P���2��ӟ����֠�[�X�8��,��اJ�#G?�~"{y����v�\���lP�;�Q8���,%���� , ��9}+D�@�6 �������A��S*R�UЉ �	����B�ͽ��Q�u�6���� �t<L� ���a���#�?̼<䓷E� y�����_FDY#o��&���	\�����$'HL�����������tJ���q�������9���F�Y�k�(������D˪~�a��J5�2
~�2�q�W���Wg`�]�c6��٘"��<��he�9��^�Lo�M���(`W͇$��@u�>��g���$��vI����Y���|���)	�4�m��p�V0��sNv��pYݲ��'��e�-�ƺ��8CK���~���l.�V(�ɕ���c��������c��U@�;�s�<��xϼ��'�j�c�ع%���g��X�L��KT��j�^�[S����%��Y&9�b�1�a}y��B.���yu��<��[���p��*�8S�K�5J�HK�+�I������=j���0�|�y}�F�3.Z��9o�
�� >.�Bm��@��`^�t
ZQ���u�����y2:�ל��{}r���Bz�'x ��7�}L#�[Z�Q_i�)�c�Iqn����x�x���9+�K�@b�^�6UK�1ǽqHfJ�( �:��`��S�5އA��b��)_H���s?�h�6�[L���z�2B�0��:����f�>������Ƿ�0��Гf�;���,�ϋ<?����& �C�7��L(�
�?�m?K��� Klp�Y�5�BX'��{ŉ7��e=��Ofйa0��>n�_�h�/�2�]��� 9��!8�$�h�ؼ�ԵV凤0�e�	t"<�)�*TG�VZ\�R���S7mw�Ex�X��������(�p<]�"T����m��WaҊ��B#�-�=]P%���X�#���#��HՋʎ�>B�+IK�̮B����\K���ҲEf�yM#abi�K��	�5Պ4#�(o��sgyӸ�ݕ���s�xO���'��F�d`cLg����	��)[W$$-�	��D�F/$�]a�ۨ���8q+��\~��i�u�)�zFv��2��9L��8DU����H������J����9 ��+_�4�BÊ>$'�1Y���3̕�~o�7F�5?�����eOx\�����k��;c"������E$� n9x�5�V��6�
�c���p��a ��ܞ�Gl͙� �����@�.�lp��H&�-L]�L���@&���ʾ�[�/^�����K�/6�f`�����z�	���F�IdY�&�Ǵ��S�A�)L=���-?j�u<�oz�["���X�dT� �{A�' �Ӑ*R�M�C����� �a��WE��/H,�4�����/Dq��\�dt��9��7�#�a���0V2�md�4�8���$ *O�x��?؝]��$�M-��'$fi���h�Ч.����g��^�3���݋P����&E�.·���l�ط�bB!4�W�Jt>eu	i�j�]��Xu8 E�k�P���ϑl�?E4h"�j4�A� \�^��T�M\Z���H��{�0��9����]�"�[���j%��x�d�q�7�����#�WTARj~/0y���"Wnr
8SQ�cW^ܫ�@�H[���?4%�ӌx��ɗ��[�Ȑ��c�	8.�p�j�� E�Ծ�z��x0�c�܂tȪL9��6ۚ�Kx�^+'\���L8���9ҳ��=|�׆Lof���R�[��~�x4 3����`�� �kHN7���s�%-ɚ�=M9E��Z!>@ s���\��ݨI
I�O��u2ú�x<e]� Tb�U�J�p�K�����.wiE�H����(bz�^Y���Mټ�R��%�n�[
9�j������z)K�;��GBEp9븐J�Js�g�Q_H���C�lhVs���~�
2af���`��D㪡-1.W�xj�UEh^�A0�Ž���c+�rS��vA/���{�	����\�#Q�\m�Fp <���_����G��!�Gb�����"��EV �m���������ȇ�7�"�٦nP�C��e{0�^�L��94�R[(U����;��$ў���2U���C��荻][,*yRM�A��a,�*��/�+$(��Gb���C1�V+l�F����F�B��"ݑh���~�;�);�
��}f������+]v�*F�+(:��Z:��O��	�R�7|�9��:���&�hq���)[�wrٳi.�H� l�(��#~ޘ,������>M�J}�ТЪ��y,��C	&�!@�GL��͠��B���v���!^X�L%�rdZ��F�bw�<�����(�~�҇�N����d�%�<��;j?�����<t�f��1�]���9G���1���r-_�`i����T�L7G&ۅ�+���}8�;BJ��R�� ��F*|=3�/�;�
��hbz�%e)���V���-��!BM�� ��=��9P�K�Ԭ�����^�^�t?�1t7B�a�Ʊ�Ѹ5�|�d�Y���ZE�%z��I�d�p/ȅ�xv��N5��+�}8�H�!���-F�y\�㞗5��0j[�ws�ܶj�,�1C��o&�>:�<E�Ed���'����%NQPC�J��ͅԊ;�d���+]}0pC+TCG�dF���߈d[��q*_F��,~�xkƸm�AftB��C��Rs� ��=�.\i�n��1J4C���]�+�x	k�YA�d��W�NDB�Ӏ����R�F� �G���K��@q�o�"�c"�7.�ͮ�$X^��I�'�&A`�"�"���+;���.U���	T������0�
�L=)��f���Zz.�~�r�3��Qi�~��Z�-ޓ�"��#�,_�QȜgS��a����O=	kfnyk�7FK��f�ָ~�q!���UF�W�Ҝ2����HS�fC`v`��������	b0��Q�V�{�C�Y� �^����}�:��^��b��g���~i)>\���Ґ� �3�/6/�'T��|�&o�~�Z�"�/��%v�?DQ�|�7Y�֗�,M���[g��&�oڌ��H0t|�y�%����_2zW�$,���tN�O,��Uo>k�[P�Yx�ic�Iơ�?���p�E>�@�]��0�0ʥ��?�<�+N[Q�!�.~�S�ܻ��{�.g5U03���n�j������)��O�/d,Ip�q6�����/��*�sO)l-{��9��܋{m�k��1D�#!�bJ�{wg�G��-L�8Қ�g<��-���%)�9C}�Y�[F|��D.�).�k��	?��1J�#8@^���\w����
n�_����.�t�۽F��q
L���B�����	U�6�`�4Ү#h���Y���5˨*��@��&�_MK��*�BŊu�c�,�DB����M�2����҄�U����i�`=�U�O�v�� '�]��պk�Д���<c�֝�}���p����FCW%~��_�������R�z>��~�	Ti;�����ￍ~�^��{���n��Y��LO�c$Z}��Z.�ɨ��ø� ˺Jrҝ96�S��!�ǂz�mmrU�9�����W�g׹걿B��d���7�ҁoE����fB��GCr�M�>�]���$���*�X}3_�#��Mݯ���xc�ȭ����E�s΢3����Vn��"�o��@b�G2�my�8	�[��v�@-<�����d��7�n�r"j�����:��f篥2\��G]����侅�m�*S�d��^�qb�7q�W��D�*�tH�
{��5����RIQ�*<UF��R�죈/����{$+��ؙǴ!��Ow(���.�-�
�E9�$������:��-{5�1@s�M��I�'����i���j�Y��zIW�F]XN�ۙ�/��K�r�lq�~�"w��
��t�I�`̓�G��LW�������5�ǾI�U)�*��E�?(�Ӛ���S<\s���N�D��9=C����Yʁ�e1a�	�S�������jD�Bz	�ӵ� ���do��Y��{AH�������ˣ�u���ݤ��h���C�_ �'3.�`���,ݟR�Έ�'�9bҘ�٤�<��k7�PL�-I�L
tpe�_�ű�;��F?�j绞�@����}�5L ���o�;�y�����ǜ��o�ߢ�cd�(��u�Un6�)2߾��v�s����Ib�x��?�h9�l.	K]`N��h�`_3�Jh���C����+$�:G�����3�Y��c� 6B��H+'׃����D���P���e;���@�XtR��oL,�����R/(\�|}�F<�1��p�/R�a�����ţ��ᥞ�+��m�$p���e�chP�=�US6�_.��~��\�Z�g��ɼ��w�S6���5���z�Ҧ*2!S�|�}�C��t�B~�$`�t�;�bU��`�.b�h���^��&�ς�c���I��eq�7��R)%�rGC�(�5�+�~�Qn��Z��[M9���B���]g�i���8R_D�W�p�9�����d���Jp�eT
(�63�[H_e����3����Z�*@��Bu:<X|s�[�Ze������^�g��[�$vf�@�W��O���#O!}~(S�HJ/(�(�@�д�*��e��3a�	����}�:�V�(�R���`��k����j��v���3��C11dQ�
_�4�(v���'){"�?�(��h50�J6倜-�<����F�;�f���Y�h,@7��X�#�-4
H����N����F�:���,¬���;���/�<��g���J��f=��B;���db����f��C��N�u� j7�&������vC��|�Cz��c���á^W8�����֎�j�(|_na�j��^��(��X: ��87#�_���'�(�fa����u�_X��ѾW��ji�s��kDGxԍ^�[)��;3�W��X%�\IZ��˒&nsv��o�v�×N�BmW���a�KP!؀3����b��W�ǳ�*ŮB6u��.U���y���i���Q��S��_��y[;���S��|�q�vmՠ�<����v�[��.��������e���&�N�d��w��9��L���Dڗ���]02\-Z
�!zX>��N���W�
��9N
O��𬶾����Z�L��F�cd�|B�:�K	���:���AܴS�4_P\c�`_W���1,&;fPp��)��֢
��+�f�6����e��> e���Ku<7qؚÚ�PyE�ͥq���=����i�,�/!Z��r4wefw�OcN�C~����|K	n�z��.Mz����@G-��H�̇�%�
e"�����j�?��ٜ�Ïf�n�E˿1�Yd�ܶA]GN�2�%��%�o͌��$6�R�J'���?LF0<����9���+yZ��X?B\� N�=��(Ykp��D����Ჹ�{8�r�#?��D�pʢ�A�{@�h?I��[EPf�,���C����d/�>���ZIs��t��8����h��X�8݉:\^xѶ�y�|�h��;�aK�c�^�I��T���i�288���_��5��Hj0��6�Q�D["���Y�X�5u7���������}��x�ԏ�?+Ȉ��겎�S�� &�����F�_�#�K������Z[*X癛��/s��_��x����.f����5J���e_V��i�t���q��lm�j�(m��x���L�_+]PyE��W�����u��d��#7��)5���mv���owN���充j��-yn*���B�3��[�q�={kE]��OD�|P�E�{ksqZ8�%���K���"��3`�4����g���L����'�g��� ��2/������{ڔjɸ�
����~�q��ET���<�:��6���{e^����z�*��������-8�.��u��qI��+�� �̋��*��gN�f�W�bC�N����}Nh�4��,� w�x�G��+������N�n�$�I��VMa�-n�#�rU)WV.@��W�;cHg_o#
��5⬚�L���V�L�a,t���%���aN�UH՘�����Ⱥ��P��%��Law�j�п�����R�mC��K��� ���$]��Y�����[��Rx>��N���f�ի�ӏ"�
c�ǪϞV3��F��_*���p0��ܾ��"�*E*=�&(J#9�$��:���z~�������+y�$&QS���sF-S���t���5�9�:��ť�_��B���+�grM�K��g��m�*vZ޴�����a�������b;��d-���NV��1�~�fB	Ḙ<��%�����7!�����?�>6{�"�1��t�i<��Jb�7<7So�`&V��F�:tdd�k�8��J/g����wl4@U�-'�����T��,����G�����/��l��^#�J�Ф�`"0���-���|�g�B���7�����rq�\魷զ������ŵ�y�"Y�n	ݲ)�����g�boA��!6��v `C�7hĊP��vʍ�
zgN���WJ�;��-UInnRJ��u������X�e=��&��M�dj,6�BΨo���p�W1�Td҅��x�o�@w�$h�򓀊{�f�Y5�NJ�x��z���A"�����Y��r�?!L��)���i����
�O�}����D�fyN��`�}�Ѥ ���e��/�}��I��!XCH��-J�*���5��d�*L%���'�&�y�I���/:"�7����i���s�8�`Y4m
S�V��ꀍ��=?5��4�͝��\�e���)��%����,nHө�q��(6gL$$��[H�{��x�d���KCߴ9|N�@�g���\?�x�����1��� ���c�u.r�ZI���{��ɒ��9m� �S��%��[qlo��Z�qD�b���O��˫�ayUݣ+�WI����1s�xt쵟���Jh�<�o3<uѝ@��5��|C%6��grk�$�^ ���=��uE��]�x���n�2�io��T�?��p�h�+�f���,.��0S�ع�e�e�x�6z�?��U��6m��ե� ZF3�2y=�I_�@�����I�X��S܅�aV�����0��kF=�o�jC�i�_Aāb4t�cǵ��9n3ȑ��~#Վ<����'v/���ۥ{o���U�d����cH�- ��;HR�Ɣ�׺��> ����/�{�O��Ba�'��;���ަ�$y�e䄠�&j����b�&W3k6~w={N@T^�y�
���-�,�ye�R�Pn+og��jȄ�1�ưs���*�5o�RjA��i��t9#��Z��!���̠`����A�*��y󡪛��� ޏ�IS!��fǀ�zO��ʹ7�q@���{�"_}<2�C	�s���� )af��-��M��V��V8�K@�N��&)唽?i6�S$����r�@h<io;-�}���ˡ+�m�VN�d
gޙGI�[�Ղ�(�A�
�><�5�5��R�u]��U��k�xm��I0���f��d�'�u7�IPv���Qɦ�l��WےS�,
m�je�Uʩ�;���><���ӹ�U��޺zD}�8�j�\��>>�n�"ᓇ�(�
s�o�E$������w�,ҕ�TtS�j�u���Ե�ܺ��E~�q����������vq����]33������OŊlJF"�[�_=ɱ*>r��p�|)�v$���P�Z�ǁ�%eW[�~�7�0�eiR�e����k��]]��;|n����V/�i
�?Q��<ÅTURT��4e���?T� �0�[T��[>�3��u]	$߰ݴ��L����(1Td�m�˲�
e��Y�����,���Э�qya�%tE��;�"�pĉ��Q�C����D��|Z�;�fL�`1���E;:-I�p@ZFW|Y�l��W�&�b�6`��g5i��OW�����p$6��J���z��=}��`A��uV,����1��HB��o�m[9- �c�"�Ќ�v��Ƶ�[�3�{4[�F�\�I�B���8�,_��'�Zg���)�޴pE�? �WDi���`�s�4���qW�qߥY(�ψx��=^D�:�
hؤ'�	m���6�=�x�Zg��edj�T��G��Ĥ)AK���(>������Y�V�G���a|����C�_��yK��"������<e &���:�
��z�36j�V1�ߏ������c4�BOʺ�X�ݧn��b����@!��|��es�ZJ�\�FZ�kw)C�>mq| ��zp��:�+�x6h�0��T�o1\i